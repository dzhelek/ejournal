ei joane
da ne se obijdame
molq te!

<3

yes


K.P
