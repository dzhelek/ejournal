yes


K.P